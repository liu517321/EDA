LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY yima IS
	PORT(A:IN STD_LOGIC;
	B:IN STD_LOGIC;
	C:IN STD_LOGIC;
	G1:IN STD_LOGIC;
	G2A:IN STD_LOGIC;
	G2B:IN STD_LOGIC;
	Y:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END yima;
	
ARCHITECTURE rtl OF yima IS
BEGIN 
	PROCESS(G1,G2A,G2B,A,B,C)
	VARIABLE COMB:STD_LOGIC_VECTOR(2 DOWNTO 0);
	BEGIN
		IF(G1='1' AND G2A='0' AND G2B='0')THEN
			COMB:=C&B&A;
			CASE COMB IS
				WHEN "000"=>Y<="11111110";
				WHEN "001"=>Y<="11111101";
				WHEN "010"=>Y<="11111011";
				WHEN "011"=>Y<="11110111";
				WHEN "100"=>Y<="11101111";
				WHEN "101"=>Y<="11011111";
				WHEN "110"=>Y<="10111111";
				WHEN "111"=>Y<="01111111";
				WHEN OTHERS=>Y<="XXXXXXXX";
			END CASE;
		ELSE
			Y<="11111111";
		END IF;
	END PROCESS;
END RTL;
